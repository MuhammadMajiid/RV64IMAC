module riscv_core_top
(
    // Global inputs
    input  wire i_riscv_core_clk,
    input  wire i_riscv_core_rst_n,
    input  wire i_riscv_core_external_interrupt,
    output wire o_riscv_core_ack,
    //Data_Cache
    output wire [63:0] o_riscv_core_dcache_raddr_axi,
    output wire [63:0] o_riscv_core_dcache_wdata,
    output wire [63:0] o_riscv_core_dcache_waddr,
    output wire o_riscv_core_dcache_raddr_valid,
    output wire o_riscv_core_dcache_wvalid,
    input  wire i_riscv_core_dcache_rready,
    input  wire i_riscv_core_dcache_wresp,
    input  wire [63:0] i_riscv_core_dcache_rdata,
    output wire [ 7 : 0] o_riscv_core_dcache_wstrb,

    //INSTR_CACHE
    output wire [63:0] o_riscv_core_icache_raddr_axi,
    output wire o_riscv_core_icache_raddr_valid,
    input  wire i_riscv_core_icache_rready,
    input  wire [63:0] i_riscv_core_icache_rdata

);

riscv_core_top_2
u_riscv_core_top_2 
(
    // Global inputs
    .i_riscv_core_clk(i_riscv_core_clk)
    ,.i_riscv_core_rst_n(i_riscv_core_rst_n)
    ,.i_riscv_core_external_interrupt(i_riscv_core_external_interrupt)
    ,.o_riscv_core_ack(o_riscv_core_ack)
    //Data_Cache
    ,.mem_read_address(o_riscv_core_dcache_raddr_axi)
    ,.o_mem_write_data(o_riscv_core_dcache_wdata)
    ,.o_mem_write_address(o_riscv_core_dcache_waddr)
    ,.mem_read_req(o_riscv_core_dcache_raddr_valid)
    ,.o_mem_write_valid(o_riscv_core_dcache_wvalid)
    ,.mem_read_done(i_riscv_core_dcache_rready)
    ,.i_mem_write_done(i_riscv_core_dcache_wresp)
    ,.i_block_from_axi_data_cache(i_riscv_core_dcache_rdata)
    ,.o_mem_write_strobe(o_riscv_core_dcache_wstrb)
  //INSTR_CACHE
    ,.o_addr_from_control_to_axi(o_riscv_core_icache_raddr_axi)
    ,.o_mem_req(o_riscv_core_icache_raddr_valid)
    ,.i_mem_done(i_riscv_core_icache_rready)
    ,.i_block_from_axi_i_cache(i_riscv_core_icache_rdata)
);
endmodule