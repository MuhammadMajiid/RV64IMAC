/*

Copyright (c) 2014-2017 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001



/*
 * AXI4-Stream UART
 */
module uart_ssh #                                                                                                           
(                                                                                                                       
    parameter block_WIDTH = 8,
    parameter CLK_RATE  = 100000000, // board internal clock (def == 100MHz)
    parameter BAUD_RATE = 115200                                                                                              
)                                                                                                                           
(                                                                                                               
    input  wire                   clk,                                                                                  
    input  wire                   rst,                                                                          

    /*                                                                                                  
     * AXI input                                                                                        
     */                                                                                         
    input  wire [block_WIDTH-1:0]  tx_data,                                         
    input  wire                   tx_valid,                                    
    output wire                   tx_ready,

    /*
     * AXI output
     */
    output wire [block_WIDTH-1:0]  rx_data,
    output wire                   rx_valid,
    input  wire                   rx_ready,

    /*
     * UART interface
     */
    input  wire                   rxd,
    output wire                   txd,

    /*
     * Status
     */
    output wire                   tx_busy,
    output wire                   rx_busy,
    output wire                   rx_overrun_error,
    output wire                   rx_frame_error

    /*
     * Configuration
     */
    //input  wire [15:0]            prescale

);
localparam prescale = CLK_RATE / BAUD_RATE;

uart_tx #(
    .block_WIDTH(block_WIDTH)
)
uart_tx_inst (
    .clk(clk),
    .rst(rst),
    // axi input
    .s_axis_tdata(tx_data),
    .s_axis_tvalid(tx_valid),
    .s_axis_tready(tx_ready),
    // output
    .txd(txd),
    // status
    .busy(tx_busy)
    // configuration
    //.prescale(prescale)
);
/*
uart_rx #(
    .block_WIDTH(block_WIDTH)
)
uart_rx_inst (
    .clk(clk),
    .rst(rst),
    // axi output
    .m_axis_tdata(rx_data),
    .m_axis_tvalid(rx_valid),
    .m_axis_tready(rx_ready),
    // input
    .rxd(rxd),
    // status
    .busy(rx_busy),
    .overrun_error(rx_overrun_error),
    .frame_error(rx_frame_error),
    // configuration
    .prescale(prescale)
);
*/
endmodule